#version 330 core
layout (location = 0) in vec2 pos;

uniform mat4 MVP;

void main()
{
	gl_Position = MVP * vec4(pos.xy, 0.0, 1.0);
}
